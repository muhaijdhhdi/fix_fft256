module fix_fft (
    input clk,
    input rstn,
    input vld_in
);

endmodule